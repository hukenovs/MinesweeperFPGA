--------------------------------------------------------------------------------
--
-- Title       : ctrl_rounds_rom
-- Design      : VGA
-- Author      : Kapitanov
-- Company     : InSys
--
-- Description : ROM generator for new rounds
--
-- Rules for ROM generator: 
--	1) 0-6 - number of mines, 7 - a mine; 8-9 - forbidden combinations
--	2) 8x8 block with "mine" or "number of mines"
--	
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity ctrl_rounds_rom is
	port(
		clk		:	in std_logic;
		addr	:	in std_logic_vector(7 downto 0);
		data	:	out std_logic_vector(23 downto 0)
	);
end ctrl_rounds_rom;

architecture ctrl_rounds_rom of ctrl_rounds_rom is

signal addr_reg	: std_logic_vector(7 downto 0);

constant N8x8	: integer:=8;
constant Ngames	: integer:=32;

type round_array_3x64xN is array (Ngames*N8x8*N8x8-1 downto 0) of integer range 0 to 7;

constant mem_init0:	round_array_3x64xN:=(
	-- game 0:
	0,0,0,0,0,0,1,7,
	0,0,0,1,1,1,2,2,
	0,0,0,1,7,2,2,7,
	0,0,0,1,2,7,2,2,
	0,1,1,1,1,1,1,0,
	0,1,7,2,7,1,1,1,
	0,1,1,2,2,2,2,7,
	0,0,0,0,1,7,2,1,
	-- game 1:
	1,1,2,7,0,0,0,0,
	1,7,3,3,2,1,0,0,
	2,3,7,2,7,1,0,0,
	7,3,2,3,1,1,0,0,
	1,2,7,2,1,1,1,0,
	0,1,1,2,7,7,1,0,
	0,0,0,1,2,2,1,0,
	0,0,0,0,0,0,0,0,
	-- game 2:
	1,1,1,1,1,1,0,0,
	1,7,1,1,7,1,0,0,
	1,1,2,2,2,1,0,0,
	0,0,1,7,1,0,0,0,
	0,1,3,3,2,0,0,0,
	0,1,7,7,2,1,1,0,
	0,2,4,4,3,7,1,0,
	0,1,7,7,2,1,1,0,
	-- game 3:
	1,1,1,0,0,1,1,1,
	1,7,2,2,1,2,7,1,
	1,2,7,2,7,3,2,1,
	0,2,2,3,2,7,1,0,
	0,1,7,2,2,1,1,0,
	1,2,3,7,1,0,0,0,
	1,7,2,1,1,0,0,0,
	1,1,1,0,0,0,0,0,
	-- game 4:
	0,0,0,0,0,0,0,0,
	0,0,1,1,1,0,0,0,
	0,1,2,7,2,1,0,0,
	1,2,7,3,7,2,1,0,
	1,7,3,4,3,7,1,0,
	1,2,7,3,7,2,1,0,
	0,1,2,7,2,1,0,0,
	0,0,1,1,1,0,0,0,
	-- game 5:
	0,2,7,2,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,3,7,3,0,0,0,0,
	0,2,7,2,0,0,0,0,
	-- game 6:
	0,0,0,0,0,0,0,0,
	0,0,1,1,1,1,1,0,
	0,0,2,7,4,7,2,0,
	0,0,3,7,6,7,3,0,
	0,0,3,7,6,7,3,0,
	0,0,2,7,4,7,2,0,
	0,0,1,2,3,2,1,0,
	0,0,0,0,0,0,0,0,	
	-- game 7:
	0,0,0,0,0,0,0,0,
	0,1,1,1,1,1,1,0,
	0,2,7,2,2,7,2,0,
	0,3,7,3,3,7,3,0,
	0,3,7,3,3,7,3,0,
	0,2,7,2,2,7,2,0,
	0,1,1,1,1,1,1,0,
	0,0,0,0,0,0,0,0,
	-- game 8:
	7,2,1,0,0,0,0,0,
	2,7,2,1,0,0,0,0,
	1,2,7,2,1,0,0,0,
	0,1,2,7,2,1,0,0,
	0,0,1,2,7,2,1,0,
	0,0,0,1,2,7,2,1,
	0,0,0,0,1,2,7,2,
	0,0,0,0,0,1,2,7,	
	-- game 9:
	0,0,0,0,0,0,0,0,
	0,1,1,1,1,1,1,0,
	0,1,7,3,3,7,1,0,
	0,1,3,7,7,3,1,0,
	0,1,3,7,7,3,1,0,
	0,1,7,3,3,7,1,0,
	0,1,1,1,1,1,1,0,
	0,0,0,0,0,0,0,0,	
	-- game A:
	1,2,1,1,0,0,0,0,
	7,2,7,1,0,0,0,0,
	2,4,2,2,0,0,0,0,
	7,2,7,1,1,1,2,1,
	1,2,1,1,1,7,2,7,
	0,0,0,0,2,2,4,2,
	0,0,0,0,1,7,2,7,
	0,0,0,0,1,1,2,1,
	-- game B:
	0,0,0,0,0,0,0,0,
	0,1,2,3,3,2,1,0,
	0,1,7,7,7,7,2,0,
	0,1,2,4,5,7,2,0,
	0,0,1,2,7,2,1,0,
	0,1,2,7,2,1,0,0,
	0,1,7,2,1,0,0,0,
	0,1,1,1,0,0,0,0,
	-- game C:
	0,0,0,0,0,1,1,1,
	0,1,1,1,1,2,7,1,
	0,1,7,2,2,7,2,1,
	0,1,2,7,3,2,1,0,
	0,1,2,3,7,2,1,0,
	1,2,7,2,2,7,1,0,
	1,7,2,1,1,1,1,0,
	1,1,1,0,0,0,0,0,	
	-- game D:
	0,0,0,0,0,0,0,0,
	0,0,1,2,3,2,1,0,
	0,0,1,7,7,7,1,0,
	0,0,1,4,7,4,1,0,
	0,0,1,4,7,4,1,0,
	0,0,1,7,7,7,1,0,
	0,0,1,2,3,2,1,0,
	0,0,0,0,0,0,0,0,
	-- game E:
	1,2,2,1,1,7,1,0,
	1,7,7,1,1,1,1,0,
	1,2,2,1,0,0,0,0,
	0,0,0,1,1,1,1,1,
	0,1,1,2,7,1,1,7,
	0,1,7,2,1,1,1,1,
	0,1,1,2,2,2,1,0,
	0,0,0,1,7,7,1,0,
	-- game F:
	1,1,1,0,0,0,0,0,
	1,7,1,0,0,0,0,0,
	3,4,3,1,0,0,0,0,
	7,7,7,1,1,2,3,2,
	2,3,2,1,1,7,7,7,
	0,0,0,0,1,3,4,3,
	0,0,0,0,0,1,7,1,
	0,0,0,0,0,1,1,1,	
	-- game 10:
	7,2,1,0,0,1,2,7,
	1,7,1,0,0,1,7,2,
	1,1,1,0,0,1,1,1,
	0,0,0,1,1,1,0,0,
	0,0,0,1,7,2,1,0,
	1,1,1,1,2,7,1,0,
	2,7,1,0,1,1,1,0,
	7,2,1,0,0,0,0,0,
	-- game 11:
	0,0,0,0,1,1,1,0,
	0,1,1,1,1,7,1,0,
	1,2,7,1,2,2,2,0,
	2,7,3,1,2,7,2,0,
	2,7,3,1,2,7,2,0,
	1,2,7,1,2,2,2,0,
	0,1,1,1,1,7,1,0,
	0,0,0,0,1,1,1,0,	
	-- game 12:
	7,1,0,0,0,1,1,1,
	1,1,0,0,0,2,7,3,
	0,0,1,1,1,2,7,7,
	0,0,1,7,1,1,2,2,
	0,1,2,2,1,0,0,0,
	0,1,7,2,0,1,1,1,
	0,1,7,2,0,1,7,1,
	0,1,1,1,0,1,1,1,
	-- game 13:
	2,7,2,1,0,0,0,0,
	7,4,7,1,0,0,0,0,
	2,7,2,1,0,0,0,0,
	1,1,1,1,1,2,1,1,
	0,0,0,1,7,3,7,1,
	0,0,0,1,3,7,2,1,
	0,0,0,1,7,2,1,0,
	0,0,0,1,1,1,0,0,
	-- game 14:
	0,0,1,1,1,1,0,0,
	0,0,1,7,7,1,0,0,
	1,1,3,4,4,3,1,1,
	1,7,2,7,7,2,7,1,
	1,1,3,4,4,3,1,1,
	0,0,1,7,7,1,0,0,
	0,0,1,1,1,1,0,0,
	0,0,0,0,0,0,0,0,	
	-- game 15:
	0,0,0,0,0,0,0,0,
	0,0,1,2,3,2,1,0,
	0,0,2,7,7,7,1,0,
	0,0,2,7,4,2,1,0,
	1,1,2,1,1,0,0,0,
	1,7,2,1,1,1,1,1,
	1,1,2,7,2,2,7,1,
	0,0,1,1,2,7,2,1,
	-- game 16:
	1,2,2,1,0,0,0,0,
	2,7,7,1,0,0,0,0,
	3,7,5,2,0,0,0,0,
	3,7,7,1,0,0,0,0,
	3,7,5,2,0,0,0,0,
	2,7,7,1,0,0,0,0,
	1,2,2,1,0,0,0,0,
	0,0,0,0,0,0,0,0,
	-- game 17:
	1,1,1,0,0,1,1,1,
	1,7,2,1,1,2,7,1,
	1,2,7,3,3,7,2,1,
	0,2,3,7,7,3,2,0,
	0,1,7,3,3,7,1,0,
	0,1,1,1,1,1,1,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	-- game 18:
	0,0,0,0,0,1,1,1,
	0,0,0,1,1,2,7,1,
	0,0,0,2,7,4,2,1,
	0,1,1,2,7,7,1,0,
	0,2,7,4,3,2,1,0,
	0,2,7,7,1,0,0,0,
	1,2,2,2,1,0,0,0,
	7,1,0,0,0,0,0,0,
	-- game 19:
	0,0,0,0,0,0,0,0,
	0,1,2,3,2,1,0,0,
	0,2,7,7,7,1,0,0,
	0,3,7,6,2,1,0,0,
	0,3,7,7,1,0,0,0,
	0,3,7,3,1,0,0,0,
	0,2,7,2,0,0,0,0,
	0,1,1,1,0,0,0,0,
	-- game 1A:
	0,0,0,0,0,0,0,0,
	0,1,1,1,1,1,1,0,
	0,1,7,1,1,7,1,0,
	0,1,2,3,3,2,1,0,
	0,0,1,7,7,1,0,0,
	0,1,2,5,5,2,1,0,
	0,1,7,7,7,7,1,0,
	0,1,2,3,3,2,1,0,
	-- game 1B:
	0,0,1,2,2,1,0,0,
	0,1,2,7,7,1,0,0,
	1,2,7,3,2,1,0,0,
	2,7,3,1,0,0,0,0,
	2,7,3,1,0,0,0,0,
	1,2,7,3,2,1,0,0,
	0,1,2,7,7,1,0,0,
	0,0,1,2,2,1,0,0,
	-- game 1C:
	0,0,0,0,0,0,0,0,
	1,2,3,2,1,0,0,0,
	1,7,7,7,4,3,2,1,
	1,2,5,7,7,7,7,1,
	0,0,2,7,4,3,2,1,
	0,0,1,1,1,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	-- game 1D:
	0,0,0,0,0,0,0,0,
	0,0,0,1,2,2,1,0,
	0,0,0,2,7,7,2,0,
	0,1,2,4,7,7,2,0,
	0,2,7,7,4,2,1,0,
	0,2,7,7,2,0,0,0,
	0,1,2,2,1,0,0,0,
	0,0,0,0,0,0,0,0,
	-- game 1E:
	7,1,0,0,0,1,1,1,
	1,1,1,1,0,1,7,1,
	1,1,7,2,1,2,1,1,
	0,1,1,2,7,2,0,0,
	0,1,1,3,7,2,0,0,
	0,1,7,3,2,1,0,0,
	0,1,2,7,1,1,1,1,
	0,0,1,1,1,1,7,1,	
	-- game 1F:
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	0,0,0,0,0,0,0,0,
	2,3,3,3,3,3,3,2,
	7,7,7,7,7,7,7,7		
	);
   
type array_3x8 		is array (N8x8-1 downto 0) of std_logic_vector(2 downto 0);
type array_3x8xN 	is array (Ngames*N8x8-1 downto 0) of array_3x8;

type array_24xN 	is array (Ngames*N8x8-1 downto 0) of std_logic_vector(23 downto 0);	
		
function read_file return array_24xN is

variable mem_inis	: round_array_3x64xN;
variable data3x8xN 	: array_3x8xN;
variable data24xN 	: array_24xN;

begin 
	mem_inis := mem_init0;
	x_loop8: for jj in 0 to Ngames*N8x8-1 loop
		for ii in 0 to N8x8-1 loop
			data3x8xN(jj)(ii) := std_logic_vector(to_unsigned(mem_init0(ii+jj*8),3));
		end loop;
	end loop;
	x_loop24: for jj in 0 to Ngames*N8x8-1 loop
		data24xN(jj) := data3x8xN(jj)(7) & data3x8xN(jj)(6) & data3x8xN(jj)(5) & data3x8xN(jj)(4) & data3x8xN(jj)(3) & data3x8xN(jj)(2) & data3x8xN(jj)(1) & data3x8xN(jj)(0);
	end loop;
	return data24xN;
end read_file;		

constant rom_data : array_24xN:=read_file;  

begin

addr_reg <= addr when rising_edge(clk);
data <= rom_data(to_integer(unsigned(addr_reg)));

end ctrl_rounds_rom;